entity PrimeDetector is
	port (SW    : in bit_vector(3 downto 0);
		  Prime : out bit);
end entity;

architecture PrimeDetector_arch of PrimeDetector is

begin

end architecture;